----------------------------------------------------------------------------------
-- Company: SCSS - Trinity College Dublin
-- Engineer: Fionn Murphy - 21363904
-- 
-- Create Date: 07.11.2022 16:03:32
-- Design Name: 
-- Module Name: DP_RippleCarryAdder32Bit_21363904_TB - Sim
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DP_RippleCarryAdder32Bit_21363904_TB is
--  Port ( ); N/A
end DP_RippleCarryAdder32Bit_21363904_TB;

architecture Sim of DP_RippleCarryAdder32Bit_21363904_TB is

--Components

    component DP_RippleCarryAdder32Bit_21363904
    port ( A : in STD_LOGIC_VECTOR (31 downto 0);
           B : in STD_LOGIC_VECTOR (31 downto 0);
           C_IN : in STD_LOGIC;
           SUM : out STD_LOGIC_VECTOR (31 downto 0);
           C_OUT : out STD_LOGIC;
           V : out STD_LOGIC);
    end component;

--Signals

    signal a_TB, b_TB : std_logic_vector (31 downto 0) := (others => '0');
    signal c_in_TB : std_logic;
    
    signal sum_TB : std_logic_vector (31 downto 0) := (others => '0');
    signal c_out_TB, v_TB : std_logic;

begin

--Unit Under Test

    uut : DP_RippleCarryAdder32Bit_21363904
    PORT MAP ( A => a_TB,
               B => b_TB,
               C_IN => c_in_TB,
               SUM => sum_TB,
               C_OUT => c_out_TB,
               V => v_TB);
    
    stim_proc : process
    begin
        
        wait for 20ns;
        --Negative + Negative with Overflow
        A_TB <= "10100000000000000000000000000000";
        B_TB <= "11000000000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Negative + Negative without Overflow
        A_TB <= "10100000000000000000000000000001";
        B_TB <= "11100000000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Positive + Positive with Overflow
        A_TB <= "00100000000000000000000000000000";
        B_TB <= "01100000000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Positive + POsitive without Overflow
        A_TB <= "00100000000000000000000000000001";
        B_TB <= "01000000000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Positive + Negative without Overflow
        A_TB <= "01000000000000000000000000000000";
        B_TB <= "11000000000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Negative + Positive without Overflow with C_IN Set
        --Worst case propogation delay
        A_TB <= "11111111111111111111111111111110";
        B_TB <= "00000000000000000000000000000001";
        C_IN_TB <= '1';
        
        wait for 360ns;
        --Student ID + Number to set C-Flag
        A_TB <= "00000001010001011111110011000000";
        B_TB <= "11111111000000000000000000000000";
        C_IN_TB <= '0';
        
        wait for 360ns;
        --Student ID + Number to set V-Flag
        A_TB <= "00000001010001011111110011000000";
        B_TB <= "01111111000000000000000000000001";
        C_IN_TB <= '0';
        
        wait for 340ns;
    
    end process;    

end Sim;
